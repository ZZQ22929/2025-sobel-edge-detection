`timescale 1ns/1ps

module tb_fifo_ctrl();

reg  sclk;
reg  rst_n;
reg  rx_flag;
reg  [7:0] rx_data;
wire area2;
wire wr_area;
wire [7:0] rgb;
wire tx_flag;
wire [7:0] tx_data;

// �ļ���ȡ����
integer input_image_file;
integer edge_result_file;
reg [7:0] image_memory [0:39999]; // 200x200����
integer i;

fifo_ctrl u_fifo_ctrl(
    .sclk(sclk),
    .rst_n(rst_n),
    .rx_flag(rx_flag),
    .rx_data(rx_data),
    .area2(area2),
    .wr_area(wr_area),
    .rgb(rgb),
    .tx_flag(tx_flag),
    .tx_data(tx_data)
);

// ʱ������ - 50MHz
initial begin
    sclk = 0;
    forever #10 sclk = ~sclk;
end

// ��ʼ��
initial begin
    rst_n = 0;
    rx_flag = 0;
    rx_data = 0;
    
    // ʹ�þ���·����ȡ����ͼ���ļ�
    $display("=== ��������ͼ�� ===");
    input_image_file = $fopen("C:/Users/HP/PycharmProjects/PythonProject7/input_image.txt", "r");
    if (input_image_file == 0) begin
        $display("����: �޷��� input_image.txt");
        $display("�����ļ�·��: C:/Users/HP/PycharmProjects/PythonProject7/input_image.txt");
        $finish;
    end
    
    // ��ȡ�������ص��ڴ�
    i = 0;
    while (!$feof(input_image_file)) begin
        if ($fscanf(input_image_file, "%d\n", image_memory[i]) == 1) begin
            i = i + 1;
            if (i % 1000 == 0) begin
                $display("�Ѷ�ȡ %0d ������...", i);
            end
        end
    end
    $fclose(input_image_file);
    $display("�ɹ����� %0d ������", i);
    
    // ��������ļ���Ҳʹ�þ���·����
    edge_result_file = $fopen("C:/Users/HP/PycharmProjects/PythonProject7/edge_result.txt", "w");
    if (edge_result_file == 0) begin
        $display("����: �޷���������ļ�");
        $finish;
    end
    
    #1000;
    rst_n = 1;
    #1000;
    
    $display("=== Sobel��Ե��⿪ʼ ===");
end

// ����������
initial begin
    // �ȴ���λ���
    #2000;
    
    // ����ͼ������
    send_image_data();
    
    #100000;
    
    $fclose(edge_result_file);
    $display("\n=== Sobel��Ե������ ===");
    $display("��Ե������ѱ��浽: C:/Users/HP/PycharmProjects/PythonProject7/edge_result.txt");
    $finish;
end

// ����ͼ����������
task send_image_data;
    integer x, y;
    begin
        $display("����ͼ�����ݵ�Sobel������...");
        
        // ����200�У�ÿ��200������
        for (y = 0; y < 200; y = y + 1) begin
            for (x = 0; x < 200; x = x + 1) begin
                rx_data = image_memory[y * 200 + x];
                rx_flag = 1;
                #20;
                rx_flag = 0;
                #80;
            end
            
            // ��ʾ����
            if (y < 5 || y % 40 == 0) begin
                $display("�Ѵ���� %0d ��", y);
            end
        end
        
        $display("ͼ�����ݷ������");
    end
endtask

// ��¼��Ե��������ļ�
always @(posedge sclk) begin
    if (u_fifo_ctrl.rd_en1) begin
        // д���Ե�����
        $fwrite(edge_result_file, "%0d\n", rgb);
    end
end

// ��ش������
reg [15:0] processed_pixels = 0;
always @(posedge sclk) begin
    if (u_fifo_ctrl.rd_en1) begin
        processed_pixels <= processed_pixels + 1;
        if (processed_pixels % 1000 == 0) begin
            $display("������ %0d ����Ե�����", processed_pixels);
        end
    end
end

endmodule