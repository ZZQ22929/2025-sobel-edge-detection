/*VGAʱ������ �� ����λ�ÿ��� �� ͼ����ʾ���� �� ��ɫ������
    ��              ��              ��            ��
ͬ���ź�       �ƶ��߼�       Sobel�����ʾ   ��̬����*/

module vga_uart(
    input   wire        sclk,
    input   wire        rst_n,
    input   wire        rx,
    output  wire        tx,
    output  wire        h_sync,
    output  wire        v_sync,
    output  wire[2:0]  r,
    output  wire[2:0]  g,
    output  wire[1:0]  b  
);
    wire        vga_clk;
    wire[7:0]   rx_data;    
    wire        po_flag;
    wire        area;
    wire[7:0]   dout;
    
    // ����FIFO�����ź�
    wire        area2;
    wire        wr_area;
    wire[7:0]   fifo_rgb;    // FIFO����ı�Ե�����

    // vga_clk��������
    vga_clk_module U1(
        .sclk(sclk),
        .rst_n(rst_n),
        .vga_clk(vga_clk)     
    );

    // vga_module��������
    vga_module U2(
        .sclk(sclk),
        .rst_n(rst_n),
        .vga_clk(vga_clk),
        .h_sync(h_sync),
        .v_sync(v_sync),
        .dout(dout),
        .r(r),
        .g(g),
        .area(area),
        .b(b)  
    );

    // uart_top��������
    uart_top U3(
        .sclk(sclk),
        .rst_n(rst_n), 
        .rx(rx),
        .tx(tx),
        .po_flag(po_flag),
        .po_data(rx_data)
    );

    // fifo_ctrl�������� - ����
    fifo_ctrl U4(
        .sclk(sclk),
        .rst_n(rst_n),
        .rx_flag(po_flag),    // ʹ��UART������ɱ�־
        .rx_data(rx_data),    // UART���յ�����
        .area2(area2),
        .wr_area(wr_area),
        .rgb(fifo_rgb)        // FIFO����ı�Ե�����
    );

    // ram_ctrl��������
    ram_ctrl U5(
        .sclk(sclk),
        .rst_n(rst_n),
        .vga_clk(vga_clk),
        .pi_flag(po_flag),
        .rgb(fifo_rgb),       // ����FIFO�����������ֱ������rx_data
        .area2(area2),
        .area(area),
        .dout(dout)
    );

endmodule