module fifo_200x8(
    input         clk,
    input  [7:0]  din,
    input         wr_en,
    input         rd_en,
    output reg [7:0]  dout,  // ��Ϊreg����
    output        full,
    output        empty
);

// FIFO����
parameter DEPTH = 200;
parameter WIDTH = 8;
parameter ADDR_WIDTH = 8;  // 2^8=256 > 200

// �ڲ��ź�
reg [WIDTH-1:0] mem [0:DEPTH-1];
reg [ADDR_WIDTH-1:0] wr_ptr = 0;
reg [ADDR_WIDTH-1:0] rd_ptr = 0;
reg [ADDR_WIDTH:0] count = 0;  // ����һλ���ڼ����/��

// д����
always @(posedge clk) begin
    if (wr_en && !full) begin
        mem[wr_ptr] <= din;
        wr_ptr <= (wr_ptr == DEPTH-1) ? 0 : wr_ptr + 1;
    end
end

// ������ - �޸���
always @(posedge clk) begin
    if (rd_en && !empty) begin
        dout <= mem[rd_ptr];
        rd_ptr <= (rd_ptr == DEPTH-1) ? 0 : rd_ptr + 1;
    end
    else if (!rd_en) begin
        // ���ֵ�ǰ���ֵ
        dout <= dout;
    end
end

// ����������
always @(posedge clk) begin
    case ({wr_en && !full, rd_en && !empty})
        2'b01: count <= count - 1;  // ֻ��
        2'b10: count <= count + 1;  // ֻд
        2'b11: count <= count;      // ͬʱ��д����������
        default: count <= count;    // �޲���
    endcase
end

// ����־
assign full = (count == DEPTH);

// �ձ�־  
assign empty = (count == 0);

endmodule