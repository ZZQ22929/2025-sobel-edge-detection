module uart_ctrl(
    input        wire        sclk,
    input        wire        rst_n,
    input        wire        rx,
    input        wire        tx_flag,    // ���� fifo_ctrl �ķ��ͱ�־
    input        wire [7:0]  tx_data,    // ���� fifo_ctrl �ķ�������
    output       wire        po_flag,
    output       wire [7:0]  rx_data,
    output       wire        tx          // TX���
);

wire                rx_bit_flag;
wire [3:0]          rx_bit_cnt;
wire                tx_bit_flag;
wire [3:0]          tx_bit_cnt;
wire                rx_flag;
wire                uart_tx_tx;  // ���� uart_tx �� tx �ź�

// bps - ��Ҫ�޸���֧��TX
uart_bps_rx U1(
    .sclk          (sclk),
    .rst_n         (rst_n),
    .rx_flag       (rx_flag),
    .tx_flag       (tx_flag),      // ʹ������ fifo_ctrl �� tx_flag
    .rx_bit_flag   (rx_bit_flag),
    .rx_bit_cnt    (rx_bit_cnt),
    .tx_bit_flag   (tx_bit_flag),
    .tx_bit_cnt    (tx_bit_cnt)
);

// rx
uart_rx U2(
    .sclk          (sclk),
    .rst_n         (rst_n),
    .rx            (rx),
    .rx_bit_cnt    (rx_bit_cnt),
    .rx_bit_flag   (rx_bit_flag),
    .po_data       (rx_data),
    .rx_flag       (rx_flag),
    .po_flag       (po_flag)
);

// tx - �޸�ʵ������ʹ������ fifo_ctrl ���ź�
uart_tx U3(
    .sclk          (sclk),
    .rst_n         (rst_n),
    .po_flag       (tx_flag),      // ʹ������ fifo_ctrl �� tx_flag ��Ϊ���ʹ���
    .po_data       (tx_data),      // ʹ������ fifo_ctrl �� tx_data
    .tx_bit_flag   (tx_bit_flag),
    .tx_bit_cnt    (tx_bit_cnt),
    .tx_flag       (),             // ���������ǲ���Ҫ
    .tx_data       (tx)            // ���ӵ��������
);

endmodule