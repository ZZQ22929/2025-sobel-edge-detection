//RX���� �� uart_rx �� �������� �� uart_tx �� TX����

module uart_top(
    input        wire        sclk,
    input        wire        rst_n, 
    input        wire        rx,
    output       wire        tx,
    output       wire        po_flag,
    output       wire[7:0]   po_data
);

// �ڲ��źŶ���
wire            rx_flag;        // ����ʹ���ź�
wire            rx_bit_flag;    // ����λ������־
wire [3:0]      rx_bit_cnt;     // ����λ������
wire            tx_flag;        // ����ʹ���ź�  
wire            tx_bit_flag;    // ����λ������־
wire [3:0]      tx_bit_cnt;     // ����λ������
wire [7:0]      rx_po_data;     // ��������

// UART����ģ��ʵ����
uart_rx u_uart_rx(
    .sclk        (sclk),
    .rst_n       (rst_n),
    .rx          (rx),
    .rx_bit_cnt  (rx_bit_cnt),
    .rx_bit_flag (rx_bit_flag),
    .po_data     (rx_po_data),
    .rx_flag     (rx_flag),
    .po_flag     (po_flag)
);

// ����������ģ��ʵ����
uart_bps_rx u_uart_bps_rx(
    .sclk        (sclk),
    .rst_n       (rst_n),
    .rx_flag     (rx_flag),
    .tx_flag     (tx_flag),
    .rx_bit_flag (rx_bit_flag),
    .rx_bit_cnt  (rx_bit_cnt),
    .tx_bit_flag (tx_bit_flag),
    .tx_bit_cnt  (tx_bit_cnt)
);

// UART����ģ��ʵ����
uart_tx u_uart_tx(
    .sclk        (sclk),
    .rst_n       (rst_n),
    .po_flag     (po_flag),        // ʹ�ý�����ɱ�־��Ϊ���ʹ���
    .po_data     (rx_po_data),     // �����յ�������ֱ�ӷ��ͻ�ȥ
    .tx_bit_flag (tx_bit_flag),
    .tx_bit_cnt  (tx_bit_cnt),
    .tx_flag     (tx_flag),
    .tx_data     (tx)
);

// ������յ�������
assign po_data = rx_po_data;

endmodule