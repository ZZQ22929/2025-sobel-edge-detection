`timescale 1ns/1ps

module tb_better_image();

reg clk, rst_n, rx;

initial begin
    clk = 0; rst_n = 0; rx = 1;
    
    $display("=== Processing Better Image ===");
    
    #1000;
    rst_n = 1;
    #1000;
    
    process_better_image();
    
    #1000;
    $display("Better image processing completed!");
    $finish;
end

task process_better_image;
    integer f_in, f_out, i;
    reg [79:0] line;
    begin
        f_in = $fopen("my_image_better.txt", "r");  // ʹ���Ż����ͼƬ
        f_out = $fopen("better_result.txt", "w");
        
        $display("Processing optimized image...");
        
        for (i = 0; i < 200; i = i + 1) begin  // �����������
            if ($fgets(line, f_in) != 0) begin
                // ģ���Ե��⣺�����شӺڱ�׻�ױ��ʱ���Ϊ��Ե
                if (i > 0) begin
                    // �򵥱�Ե����߼�
                    if (line[1:0] == "FF") 
                        $fdisplay(f_out, "FF");  // ��ɫ����
                    else
                        $fdisplay(f_out, "00");  // ��ɫ����
                end
                
                if (i % 40 == 0)
                    $display("  Processed %d/200 pixels", i);
            end
        end
        
        $fclose(f_in);
        $fclose(f_out);
        $display("Generated: better_result.txt");
    end
endtask

always #10 clk = ~clk;

endmodule