`timescale 1ns/1ps

module tb_vga_uart();

reg  sclk;
reg  rst_n;
reg  rx;
wire tx;
wire h_sync;
wire v_sync;
wire [2:0] r;
wire [2:0] g;
wire [1:0] b;

// ���ڼ���źű��صļĴ���
reg h_sync_prev;
reg v_sync_prev;

vga_uart u_vga_uart(
    .sclk(sclk),
    .rst_n(rst_n),
    .rx(rx),
    .tx(tx),
    .h_sync(h_sync),
    .v_sync(v_sync),
    .r(r),
    .g(g),
    .b(b)
);

// ϵͳʱ�� 50MHz
initial begin
    sclk = 0;
    forever #10 sclk = ~sclk;
end

// ��ʼ��
initial begin
    rst_n = 0;
    rx = 1;
    h_sync_prev = 0;
    v_sync_prev = 0;
    #1000;
    rst_n = 1;
    #1000;
    
    $display("=== VGA UART System Test Start ===");
    $display("Time: %0t ns", $time);
end

// ����������
initial begin
    // �ȴ���λ���
    #2000;
    
    // ���ԣ�����200x200ͼ�����ϵͳ
    $display("\n--- Test: 200x200 Image Transmission ---");
    test_large_image();
    
    #1000000;  // �ӳ�����ʱ��۲�VGA���
    
    $display("\n=== VGA UART System Test Completed ===");
    $display("Time: %0t ns", $time);
    $finish;
end

// ���ʹ�ͼ�����
task test_large_image;
    integer i, j;
    begin
        $display("Sending 200x200 test image via UART...");
        
        // ����200x200����ͼ��
        for (j = 0; j < 200; j = j + 1) begin
            for (i = 0; i < 200; i = i + 1) begin
                // �������Եı�Ե����ͼ��
                if (i < 100)  // ��벿�ֺ�ɫ���Ұ벿�ְ�ɫ��������ֱ��Ե
                    send_byte(8'h00);  // ��ɫ
                else
                    send_byte(8'hFF);  // ��ɫ
                
                #500;  // �ֽڼ���
            end
            if (j % 20 == 0) begin
                $display("  Line %0d sent", j);
            end
        end
        
        $display("Large image transmission completed");
    end
endtask

// ���͵����ֽ�
task send_byte;
    input [7:0] data;
    integer k;
    begin
        // ��ʼλ
        rx = 1'b0;
        #8680;
        
        // 8������λ (LSB first)
        for (k = 0; k < 8; k = k + 1) begin
            rx = data[k];
            #8680;
        end
        
        // ֹͣλ
        rx = 1'b1;
        #8680;
    end
endtask

// ����źű���
always @(posedge sclk) begin
    h_sync_prev <= h_sync;
    v_sync_prev <= v_sync;
    
    // ��ʾVGAͬ���źű仯
    if (h_sync && !h_sync_prev) begin
        $display("H_SYNC: rising edge");
    end
    if (v_sync && !v_sync_prev) begin
        $display("V_SYNC: rising edge - FRAME START");
    end
end

// ���RGB��� - ֻ���б仯ʱ��ʾ
reg [7:0] last_rgb;
always @(posedge sclk) begin
    last_rgb <= {r, g, b};
    if ({r, g, b} !== last_rgb && (r != 0 || g != 0 || b != 0)) begin
        $display("RGB_CHANGE: r=%b, g=%b, b=%b", r, g, b);
    end
end

// ���ϵͳ״̬
always @(posedge sclk) begin
    // ��ʾUART����
    if (u_vga_uart.U3.po_flag) begin
        $display("UART_RX: data=0x%h", u_vga_uart.U3.po_data);
    end
end

// ���α���
initial begin
    $dumpfile("vga_uart.vcd");
    $dumpvars(0, tb_vga_uart);
end

endmodule