/*����ʱ����(sclk) �� ˫�˿�RAM �� ��ʾʱ����(vga_clk)
     ��                    ��              ��
 Sobel������ �� ֡���� �� VGA��ʾ����*/

module ram_39204x8(
    input         clka,
    input         wea,
    input  [15:0] addra,
    input  [7:0]  dina,
    input         clkb,
    input  [15:0] addrb,
    output reg [7:0] doutb
);

// RAM����
parameter DEPTH = 39204;
parameter WIDTH = 8;
parameter ADDR_WIDTH = 16;

// RAM�洢��
reg [WIDTH-1:0] mem [0:DEPTH-1];

// д���� (�˿�A)
always @(posedge clka) begin
    if (wea) begin
        if (addra < DEPTH) begin
            mem[addra] <= dina;
        end
    end
end

// ������ (�˿�B)
always @(posedge clkb) begin
    if (addrb < DEPTH) begin
        doutb <= mem[addrb];
    end else begin
        doutb <= 8'h00;  // ��ַԽ��ʱ���0
    end
end

endmodule